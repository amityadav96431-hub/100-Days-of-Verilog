module not_gate_behavioral(
  input a,
  output y
);
  assign y = ~a;
endmodule
